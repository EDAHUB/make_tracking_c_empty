// DESCRIPTION: Verilator: Verilog Test module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2003 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0
// ======================================================================

module sub
  (
   input clk /*verilator public*/,
   input reset_l/*verilator public*/,
   input  [31:0] in_small/*verilator public*/,
   output [31:0] out_small/*verilator public*/
   );


endmodule
